library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity VGA  is

	port(	clk  		: in std_logic;
			scoreVGA	: in	integer;
			quadrante: in std_logic_vector(3 downto 0);
			red   	: out std_logic_vector(2 downto 0);
			green 	: out std_logic_vector(2 downto 0);
			blue  	: out std_logic_vector(1 downto 0);
			hs    	: out std_logic;
			vs    	: out std_logic
			);
end VGA ;
-- gerenciamento das rotinas para comunica��o com monitor (VGA)
architecture Behavioral of VGA is
	-- criando "tipo" para matriz binaria que gera a imagem do n�mero
	type valor is array (0 to 97) of std_logic_vector (0 to 63);
	
	-- constante para matriz do n�mero 0
	constant valor0 : valor := (
	"0000000000000000000000000011111111111100000000000000000000000000",
	"0000000000000000000000111111111111111111110000000000000000000000",
	"0000000000000000000011111111111111111111111100000000000000000000",
	"0000000000000000001111111111111111111111111111000000000000000000",
	"0000000000000000111111111111111111111111111111110000000000000000",
	"0000000000000001111111111111111111111111111111111000000000000000",
	"0000000000000111111111111111111111111111111111111100000000000000",
	"0000000000001111111111111111111111111111111111111111000000000000",
	"0000000000011111111111111111111111111111111111111111000000000000",
	"0000000000011111111111111111111111111111111111111111100000000000",
	"0000000000111111111111111111111111111111111111111111110000000000",
	"0000000001111111111111111111111111111111111111111111111000000000",
	"0000000001111111111111111111111111111111111111111111111000000000",
	"0000000011111111111111111111111111111111111111111111111100000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000001111111111111111111111100000011111111111111111111111000000",
	"0000001111111111111111111110000000000111111111111111111111000000",
	"0000001111111111111111111100000000000011111111111111111111000000",
	"0000011111111111111111111000000000000001111111111111111111100000",
	"0000011111111111111111110000000000000000111111111111111111100000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000111111111111111111000000000000000000001111111111111111110000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111110000000000000000000000111111111111111111000",
	"0001111111111111111110000000000000000000000111111111111111111000",
	"0001111111111111111110000000000000000000000111111111111111111000",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000011111111111111111100",
	"0011111111111111111100000000000000000000000011111111111111111100",
	"0011111111111111111100000000000000000000000011111111111111111100",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0011111111111111111100000000000000000000000011111111111111111100",
	"0011111111111111111100000000000000000000000011111111111111111100",
	"0011111111111111111100000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111000",
	"0001111111111111111110000000000000000000000111111111111111111000",
	"0001111111111111111110000000000000000000000111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111110000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000011111111111111111110000000000000000111111111111111111100000",
	"0000011111111111111111111000000000000001111111111111111111100000",
	"0000011111111111111111111100000000000011111111111111111111000000",
	"0000001111111111111111111110000000000111111111111111111111000000",
	"0000001111111111111111111111100000011111111111111111111111000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000000011111111111111111111111111111111111111111111111100000000",
	"0000000011111111111111111111111111111111111111111111111000000000",
	"0000000001111111111111111111111111111111111111111111111000000000",
	"0000000000111111111111111111111111111111111111111111110000000000",
	"0000000000011111111111111111111111111111111111111111100000000000",
	"0000000000001111111111111111111111111111111111111111100000000000",
	"0000000000000111111111111111111111111111111111111111000000000000",
	"0000000000000011111111111111111111111111111111111110000000000000",
	"0000000000000001111111111111111111111111111111111000000000000000",
	"0000000000000000111111111111111111111111111111110000000000000000",
	"0000000000000000001111111111111111111111111111000000000000000000",
	"0000000000000000000011111111111111111111111100000000000000000000",
	"0000000000000000000000111111111111111111110000000000000000000000",
	"0000000000000000000000000011111111111100000000000000000000000000");
	
	-- constante para matriz do n�mero 1
	constant valor1 : valor := (
	"0000000000000000000000000000111111111111111000000000000000000000",
	"0000000000000000000000000000111111111111111000000000000000000000",
	"0000000000000000000000000001111111111111111000000000000000000000",
	"0000000000000000000000000001111111111111111000000000000000000000",
	"0000000000000000000000000011111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000001111111111111111111000000000000000000000",
	"0000000000000000000000011111111111111111111000000000000000000000",
	"0000000000000000000000011111111111111111111000000000000000000000",
	"0000000000000000000000111111111111111111111000000000000000000000",
	"0000000000000000000001111111111111111111111000000000000000000000",
	"0000000000000000000011111111111111111111111000000000000000000000",
	"0000000000000000000111111111111111111111111000000000000000000000",
	"0000000000000000011111111111111111111111111000000000000000000000",
	"0000000000000000111111111111111111111111111000000000000000000000",
	"0000000000000001111111111111111111111111111000000000000000000000",
	"0000000000000111111111111111111111111111111000000000000000000000",
	"0000000000001111111111111111111111111111111000000000000000000000",
	"0000000000111111111111111111111111111111111000000000000000000000",
	"0000000001111111111111111111111111111111111000000000000000000000",
	"0000000111111111111111111111111111111111111000000000000000000000",
	"0000011111111111111111111111111111111111111000000000000000000000",
	"0011111111111111111111111111111111111111111000000000000000000000",
	"0111111111111111111111111111111111111111111000000000000000000000",
	"0111111111111111111111111111111111111111111000000000000000000000",
	"0111111111111111111111111111111111111111111000000000000000000000",
	"0111111111111111111111110111111111111111111000000000000000000000",
	"0111111111111111111111100111111111111111111000000000000000000000",
	"0111111111111111111111000111111111111111111000000000000000000000",
	"0111111111111111111110000111111111111111111000000000000000000000",
	"0111111111111111111100000111111111111111111000000000000000000000",
	"0111111111111111111000000111111111111111111000000000000000000000",
	"0111111111111111100000000111111111111111111000000000000000000000",
	"0111111111111111000000000111111111111111111000000000000000000000",
	"0111111111111100000000000111111111111111111000000000000000000000",
	"0111111111111000000000000111111111111111111000000000000000000000",
	"0111111111100000000000000111111111111111111000000000000000000000",
	"0111111110000000000000000111111111111111111000000000000000000000",
	"0111111000000000000000000111111111111111111000000000000000000000",
	"0111100000000000000000000111111111111111111000000000000000000000",
	"0100000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111111000000000000000000000",
	"0000000000000000000000000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000000000000000000000000");
	
	-- constante para matriz do n�mero 2
	constant valor2 : valor := (
	"0000000000000000000000000001111111111111000000000000000000000000",
	"0000000000000000000000011111111111111111111110000000000000000000",
	"0000000000000000000011111111111111111111111111110000000000000000",
	"0000000000000000001111111111111111111111111111111100000000000000",
	"0000000000000000111111111111111111111111111111111110000000000000",
	"0000000000000011111111111111111111111111111111111111100000000000",
	"0000000000000111111111111111111111111111111111111111110000000000",
	"0000000000001111111111111111111111111111111111111111111000000000",
	"0000000000011111111111111111111111111111111111111111111100000000",
	"0000000000111111111111111111111111111111111111111111111110000000",
	"0000000001111111111111111111111111111111111111111111111111000000",
	"0000000011111111111111111111111111111111111111111111111111100000",
	"0000000011111111111111111111111111111111111111111111111111100000",
	"0000000111111111111111111111111111111111111111111111111111110000",
	"0000000111111111111111111111111111111111111111111111111111110000",
	"0000001111111111111111111111111111111111111111111111111111111000",
	"0000001111111111111111111111110000000111111111111111111111111000",
	"0000011111111111111111111110000000000001111111111111111111111100",
	"0000011111111111111111111100000000000000111111111111111111111100",
	"0000011111111111111111111000000000000000011111111111111111111100",
	"0000111111111111111111110000000000000000001111111111111111111100",
	"0000111111111111111111110000000000000000000111111111111111111110",
	"0000111111111111111111100000000000000000000111111111111111111110",
	"0000111111111111111111100000000000000000000111111111111111111110",
	"0000111111111111111111100000000000000000000011111111111111111110",
	"0001111111111111111111100000000000000000000011111111111111111110",
	"0001111111111111111111000000000000000000000011111111111111111110",
	"0001111111111111111111000000000000000000000011111111111111111110",
	"0000011111111111111111000000000000000000000011111111111111111110",
	"0000000000000000111111000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111100",
	"0000000000000000000000000000000000000000000111111111111111111100",
	"0000000000000000000000000000000000000000000111111111111111111100",
	"0000000000000000000000000000000000000000000111111111111111111100",
	"0000000000000000000000000000000000000000001111111111111111111000",
	"0000000000000000000000000000000000000000001111111111111111111000",
	"0000000000000000000000000000000000000000011111111111111111111000",
	"0000000000000000000000000000000000000000011111111111111111110000",
	"0000000000000000000000000000000000000000111111111111111111110000",
	"0000000000000000000000000000000000000001111111111111111111100000",
	"0000000000000000000000000000000000000011111111111111111111100000",
	"0000000000000000000000000000000000000111111111111111111111000000",
	"0000000000000000000000000000000000000111111111111111111111000000",
	"0000000000000000000000000000000000001111111111111111111110000000",
	"0000000000000000000000000000000000011111111111111111111110000000",
	"0000000000000000000000000000000000111111111111111111111100000000",
	"0000000000000000000000000000000001111111111111111111111000000000",
	"0000000000000000000000000000000011111111111111111111111000000000",
	"0000000000000000000000000000000111111111111111111111110000000000",
	"0000000000000000000000000000001111111111111111111111100000000000",
	"0000000000000000000000000000011111111111111111111111000000000000",
	"0000000000000000000000000000111111111111111111111110000000000000",
	"0000000000000000000000000001111111111111111111111110000000000000",
	"0000000000000000000000000011111111111111111111111100000000000000",
	"0000000000000000000000000111111111111111111111111000000000000000",
	"0000000000000000000000001111111111111111111111110000000000000000",
	"0000000000000000000000011111111111111111111111100000000000000000",
	"0000000000000000000000111111111111111111111111000000000000000000",
	"0000000000000000000001111111111111111111111110000000000000000000",
	"0000000000000000000011111111111111111111111000000000000000000000",
	"0000000000000000000111111111111111111111110000000000000000000000",
	"0000000000000000001111111111111111111111100000000000000000000000",
	"0000000000000000011111111111111111111111000000000000000000000000",
	"0000000000000000111111111111111111111110000000000000000000000000",
	"0000000000000001111111111111111111111100000000000000000000000000",
	"0000000000000001111111111111111111111000000000000000000000000000",
	"0000000000000011111111111111111111110000000000000000000000000000",
	"0000000000000111111111111111111111100000000000000000000000000000",
	"0000000000001111111111111111111111000000000000000000000000000000",
	"0000000000011111111111111111111110000000000000000000000000000000",
	"0000000000111111111111111111111100000000000000000000000000000000",
	"0000000000111111111111111111111000000000000000000000000000000000",
	"0000000001111111111111111111111000000000000000000000000000000000",
	"0000000011111111111111111111110000000000000000000000000000000000",
	"0000000011111111111111111111100000000000000000000000000000000000",
	"0000000111111111111111111111100000000000000000000000000000000000",
	"0000000111111111111111111111111111111111111111111111111111111110",
	"0000001111111111111111111111111111111111111111111111111111111110",
	"0000011111111111111111111111111111111111111111111111111111111110",
	"0000011111111111111111111111111111111111111111111111111111111110",
	"0000011111111111111111111111111111111111111111111111111111111110",
	"0000111111111111111111111111111111111111111111111111111111111110",
	"0000111111111111111111111111111111111111111111111111111111111110",
	"0001111111111111111111111111111111111111111111111111111111111110",
	"0001111111111111111111111111111111111111111111111111111111111110",
	"0001111111111111111111111111111111111111111111111111111111111110",
	"0011111111111111111111111111111111111111111111111111111111111110",
	"0011111111111111111111111111111111111111111111111111111111111110",
	"0011111111111111111111111111111111111111111111111111111111111110",
	"0011111111111111111111111111111111111111111111111111111111111110",
	"0011111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110");
	
	-- constante para matriz do n�mero 3
	constant valor3 : valor := (
	"0000000000000000000000000011111111111100000000000000000000000000",
	"0000000000000000000001111111111111111111110000000000000000000000",
	"0000000000000000000111111111111111111111111100000000000000000000",
	"0000000000000000011111111111111111111111111111000000000000000000",
	"0000000000000001111111111111111111111111111111110000000000000000",
	"0000000000000011111111111111111111111111111111111000000000000000",
	"0000000000001111111111111111111111111111111111111100000000000000",
	"0000000000011111111111111111111111111111111111111110000000000000",
	"0000000000111111111111111111111111111111111111111111000000000000",
	"0000000001111111111111111111111111111111111111111111100000000000",
	"0000000001111111111111111111111111111111111111111111110000000000",
	"0000000011111111111111111111111111111111111111111111111000000000",
	"0000000111111111111111111111111111111111111111111111111000000000",
	"0000000111111111111111111111111111111111111111111111111100000000",
	"0000001111111111111111111111111111111111111111111111111110000000",
	"0000001111111111111111111111111111111111111111111111111110000000",
	"0000011111111111111111111111100000011111111111111111111110000000",
	"0000011111111111111111111110000000001111111111111111111111000000",
	"0000011111111111111111111100000000000011111111111111111111000000",
	"0000111111111111111111111000000000000011111111111111111111000000",
	"0000111111111111111111110000000000000001111111111111111111100000",
	"0000111111111111111111110000000000000001111111111111111111100000",
	"0000111111111111111111100000000000000000111111111111111111100000",
	"0001111111111111111111100000000000000000111111111111111111100000",
	"0001111111111111111111100000000000000000111111111111111111100000",
	"0000111111111111111111000000000000000000111111111111111111100000",
	"0000000000011111111111000000000000000000111111111111111111100000",
	"0000000000000000001111000000000000000000111111111111111111100000",
	"0000000000000000000000000000000000000000111111111111111111100000",
	"0000000000000000000000000000000000000000111111111111111111000000",
	"0000000000000000000000000000000000000001111111111111111111000000",
	"0000000000000000000000000000000000000001111111111111111111000000",
	"0000000000000000000000000000000000000001111111111111111110000000",
	"0000000000000000000000000000000000000011111111111111111110000000",
	"0000000000000000000000000000000000000111111111111111111100000000",
	"0000000000000000000000000000000000001111111111111111111100000000",
	"0000000000000000000000000000000000011111111111111111111000000000",
	"0000000000000000000000000000000011111111111111111111110000000000",
	"0000000000000000000000000000111111111111111111111111100000000000",
	"0000000000000000000000000001111111111111111111111111000000000000",
	"0000000000000000000000000001111111111111111111111110000000000000",
	"0000000000000000000000000001111111111111111111111100000000000000",
	"0000000000000000000000000001111111111111111111111000000000000000",
	"0000000000000000000000000001111111111111111111100000000000000000",
	"0000000000000000000000000001111111111111111110000000000000000000",
	"0000000000000000000000000001111111111111111111100000000000000000",
	"0000000000000000000000000001111111111111111111111100000000000000",
	"0000000000000000000000000001111111111111111111111111000000000000",
	"0000000000000000000000000001111111111111111111111111100000000000",
	"0000000000000000000000000011111111111111111111111111111000000000",
	"0000000000000000000000000011111111111111111111111111111100000000",
	"0000000000000000000000000011111111111111111111111111111110000000",
	"0000000000000000000000000011100000001111111111111111111111000000",
	"0000000000000000000000000000000000000011111111111111111111100000",
	"0000000000000000000000000000000000000000111111111111111111100000",
	"0000000000000000000000000000000000000000111111111111111111110000",
	"0000000000000000000000000000000000000000011111111111111111110000",
	"0000000000000000000000000000000000000000001111111111111111111000",
	"0000000000000000000000000000000000000000001111111111111111111000",
	"0000000000000000000000000000000000000000000111111111111111111100",
	"0000000000000000000000000000000000000000000111111111111111111100",
	"0000000000000000000000000000000000000000000111111111111111111100",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000111100000000000000000000000011111111111111111110",
	"0000000111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111110000000000000000000000011111111111111111110",
	"0111111111111111111110000000000000000000000111111111111111111110",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111111000000000000000000000111111111111111111100",
	"0011111111111111111111000000000000000000001111111111111111111100",
	"0011111111111111111111100000000000000000001111111111111111111100",
	"0001111111111111111111100000000000000000011111111111111111111000",
	"0001111111111111111111110000000000000000111111111111111111111000",
	"0001111111111111111111111000000000000001111111111111111111111000",
	"0000111111111111111111111110000000000011111111111111111111110000",
	"0000111111111111111111111111100000011111111111111111111111110000",
	"0000011111111111111111111111111111111111111111111111111111100000",
	"0000011111111111111111111111111111111111111111111111111111100000",
	"0000001111111111111111111111111111111111111111111111111111000000",
	"0000001111111111111111111111111111111111111111111111111110000000",
	"0000000111111111111111111111111111111111111111111111111100000000",
	"0000000011111111111111111111111111111111111111111111111100000000",
	"0000000001111111111111111111111111111111111111111111111000000000",
	"0000000000111111111111111111111111111111111111111111110000000000",
	"0000000000011111111111111111111111111111111111111111100000000000",
	"0000000000001111111111111111111111111111111111111110000000000000",
	"0000000000000111111111111111111111111111111111111100000000000000",
	"0000000000000001111111111111111111111111111111110000000000000000",
	"0000000000000000011111111111111111111111111111100000000000000000",
	"0000000000000000000111111111111111111111111110000000000000000000",
	"0000000000000000000001111111111111111111110000000000000000000000",
	"0000000000000000000000000011111111111100000000000000000000000000");
	
	-- constante para matriz do n�mero 4
	constant valor4 : valor := (
	"0000000000000000000000000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000111111111111111100000000",
	"0000000000000000000000000000000000000001111111111111111100000000",
	"0000000000000000000000000000000000000001111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000111111111111111111100000000",
	"0000000000000000000000000000000000000111111111111111111100000000",
	"0000000000000000000000000000000000001111111111111111111100000000",
	"0000000000000000000000000000000000011111111111111111111100000000",
	"0000000000000000000000000000000000011111111111111111111100000000",
	"0000000000000000000000000000000000111111111111111111111100000000",
	"0000000000000000000000000000000001111111111111111111111100000000",
	"0000000000000000000000000000000001111111111111111111111100000000",
	"0000000000000000000000000000000011111111111111111111111100000000",
	"0000000000000000000000000000000111111111111111111111111100000000",
	"0000000000000000000000000000001111111111111111111111111100000000",
	"0000000000000000000000000000001111111111111111111111111100000000",
	"0000000000000000000000000000011111111111111111111111111100000000",
	"0000000000000000000000000000111111111111111111111111111100000000",
	"0000000000000000000000000000111111111111111111111111111100000000",
	"0000000000000000000000000001111111111111111111111111111100000000",
	"0000000000000000000000000011111111111111111111111111111100000000",
	"0000000000000000000000000011111111111111111111111111111100000000",
	"0000000000000000000000000111111111111111111111111111111100000000",
	"0000000000000000000000001111111111111111111111111111111100000000",
	"0000000000000000000000001111111111111111111111111111111100000000",
	"0000000000000000000000011111111111111111111111111111111100000000",
	"0000000000000000000000111111111111111111111111111111111100000000",
	"0000000000000000000000111111111111111111111111111111111100000000",
	"0000000000000000000001111111111111111111111111111111111100000000",
	"0000000000000000000011111111111111111011111111111111111100000000",
	"0000000000000000000011111111111111110011111111111111111100000000",
	"0000000000000000000111111111111111110011111111111111111100000000",
	"0000000000000000001111111111111111100011111111111111111100000000",
	"0000000000000000011111111111111111000011111111111111111100000000",
	"0000000000000000011111111111111111000011111111111111111100000000",
	"0000000000000000111111111111111110000011111111111111111100000000",
	"0000000000000001111111111111111100000011111111111111111100000000",
	"0000000000000001111111111111111000000011111111111111111100000000",
	"0000000000000011111111111111111000000011111111111111111100000000",
	"0000000000000111111111111111110000000011111111111111111100000000",
	"0000000000000111111111111111100000000011111111111111111100000000",
	"0000000000001111111111111111100000000011111111111111111100000000",
	"0000000000011111111111111111000000000011111111111111111100000000",
	"0000000000011111111111111110000000000011111111111111111100000000",
	"0000000000111111111111111110000000000011111111111111111100000000",
	"0000000001111111111111111100000000000011111111111111111100000000",
	"0000000001111111111111111000000000000011111111111111111100000000",
	"0000000011111111111111111000000000000011111111111111111100000000",
	"0000000111111111111111110000000000000011111111111111111100000000",
	"0000000111111111111111100000000000000011111111111111111100000000",
	"0000001111111111111111100000000000000011111111111111111100000000",
	"0000011111111111111111000000000000000011111111111111111100000000",
	"0000111111111111111110000000000000000011111111111111111100000000",
	"0000111111111111111110000000000000000011111111111111111100000000",
	"0001111111111111111100000000000000000011111111111111111100000000",
	"0011111111111111111000000000000000000011111111111111111100000000",
	"0011111111111111110000000000000000000011111111111111111100000000",
	"0111111111111111110000000000000000000011111111111111111100000000",
	"1111111111111111100000000000000000000011111111111111111100000000",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000000000000000000000000");
	
	-- constante para matriz do n�mero 5
	constant valor5 : valor := (
	"0000000000000000000000000000000000000000000000000000000000000000",
	"0000000000000111111111111111111111111111111111111111111111110000",
	"0000000000000111111111111111111111111111111111111111111111110000",
	"0000000000001111111111111111111111111111111111111111111111110000",
	"0000000000001111111111111111111111111111111111111111111111110000",
	"0000000000001111111111111111111111111111111111111111111111110000",
	"0000000000001111111111111111111111111111111111111111111111110000",
	"0000000000001111111111111111111111111111111111111111111111110000",
	"0000000000011111111111111111111111111111111111111111111111110000",
	"0000000000011111111111111111111111111111111111111111111111110000",
	"0000000000011111111111111111111111111111111111111111111111110000",
	"0000000000011111111111111111111111111111111111111111111111110000",
	"0000000000011111111111111111111111111111111111111111111111110000",
	"0000000000111111111111111111111111111111111111111111111111110000",
	"0000000000111111111111111111111111111111111111111111111111110000",
	"0000000000111111111111111111111111111111111111111111111111110000",
	"0000000000111111111111111111111111111111111111111111111111110000",
	"0000000000111111111111111111111111111111111111111111111111110000",
	"0000000001111111111111111111111111111111111111111111111111110000",
	"0000000001111111111111111111111111111111111111111111111111110000",
	"0000000001111111111111111111000000000000000000000000000000000000",
	"0000000001111111111111111111000000000000000000000000000000000000",
	"0000000001111111111111111111000000000000000000000000000000000000",
	"0000000011111111111111111110000000000000000000000000000000000000",
	"0000000011111111111111111110000000000000000000000000000000000000",
	"0000000011111111111111111110000000000000000000000000000000000000",
	"0000000011111111111111111110000000000000000000000000000000000000",
	"0000000111111111111111111110000000000000000000000000000000000000",
	"0000000111111111111111111100000000000000000000000000000000000000",
	"0000000111111111111111111100000000000000000000000000000000000000",
	"0000000111111111111111111100000000000000000000000000000000000000",
	"0000000111111111111111111100000000000000000000000000000000000000",
	"0000001111111111111111111000000000000000000000000000000000000000",
	"0000001111111111111111111000000011111111110000000000000000000000",
	"0000001111111111111111111000011111111111111110000000000000000000",
	"0000001111111111111111111011111111111111111111110000000000000000",
	"0000001111111111111111111111111111111111111111111100000000000000",
	"0000011111111111111111111111111111111111111111111110000000000000",
	"0000011111111111111111111111111111111111111111111111100000000000",
	"0000011111111111111111111111111111111111111111111111110000000000",
	"0000011111111111111111111111111111111111111111111111111000000000",
	"0000011111111111111111111111111111111111111111111111111100000000",
	"0000111111111111111111111111111111111111111111111111111110000000",
	"0000111111111111111111111111111111111111111111111111111111000000",
	"0000111111111111111111111111111111111111111111111111111111000000",
	"0000111111111111111111111111111111111111111111111111111111100000",
	"0000111111111111111111111111111111111111111111111111111111110000",
	"0001111111111111111111111111111111111111111111111111111111110000",
	"0001111111111111111111111111111111111111111111111111111111111000",
	"0001111111111111111111111111000000001111111111111111111111111000",
	"0001111111111111111111111000000000000011111111111111111111111100",
	"0011111111111111111111100000000000000000111111111111111111111100",
	"0011111111111111111111000000000000000000011111111111111111111100",
	"0011111111111111111110000000000000000000001111111111111111111110",
	"0000000111111111111100000000000000000000000111111111111111111110",
	"0000000000000001111000000000000000000000000111111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111111",
	"0000000000000000000000000000000000000000000001111111111111111111",
	"0000000000000000000000000000000000000000000001111111111111111111",
	"0000000000000000000000000000000000000000000001111111111111111111",
	"0000000000000000000000000000000000000000000001111111111111111111",
	"0000000000000000000000000000000000000000000001111111111111111111",
	"0000000000000000000000000000000000000000000001111111111111111111",
	"0000000000000000000000000000000000000000000001111111111111111111",
	"0000000000000000000000000000000000000000000001111111111111111111",
	"0000000000001111000000000000000000000000000001111111111111111111",
	"0000111111111111000000000000000000000000000001111111111111111111",
	"1111111111111111000000000000000000000000000001111111111111111111",
	"1111111111111111100000000000000000000000000011111111111111111110",
	"1111111111111111100000000000000000000000000011111111111111111110",
	"0111111111111111110000000000000000000000000011111111111111111110",
	"0111111111111111110000000000000000000000000111111111111111111110",
	"0111111111111111111000000000000000000000000111111111111111111100",
	"0111111111111111111000000000000000000000001111111111111111111100",
	"0011111111111111111100000000000000000000011111111111111111111100",
	"0011111111111111111110000000000000000000111111111111111111111000",
	"0011111111111111111111100000000000000001111111111111111111111000",
	"0001111111111111111111110000000000000111111111111111111111110000",
	"0001111111111111111111111110000000111111111111111111111111110000",
	"0000111111111111111111111111111111111111111111111111111111100000",
	"0000111111111111111111111111111111111111111111111111111111100000",
	"0000011111111111111111111111111111111111111111111111111111000000",
	"0000001111111111111111111111111111111111111111111111111110000000",
	"0000001111111111111111111111111111111111111111111111111110000000",
	"0000000111111111111111111111111111111111111111111111111100000000",
	"0000000011111111111111111111111111111111111111111111111000000000",
	"0000000001111111111111111111111111111111111111111111110000000000",
	"0000000000111111111111111111111111111111111111111111100000000000",
	"0000000000011111111111111111111111111111111111111111000000000000",
	"0000000000000111111111111111111111111111111111111100000000000000",
	"0000000000000011111111111111111111111111111111111000000000000000",
	"0000000000000000111111111111111111111111111111100000000000000000",
	"0000000000000000001111111111111111111111111110000000000000000000",
	"0000000000000000000001111111111111111111110000000000000000000000",
	"0000000000000000000000000111111111111100000000000000000000000000",
	"0000000000000000000000000000000000000000000000000000000000000000");
	
	-- constante para matriz do n�mero 6
	constant valor6 : valor := (
	"0000000000000000000000000000111111111110000000000000000000000000",
	"0000000000000000000000001111111111111111111000000000000000000000",
	"0000000000000000000001111111111111111111111111000000000000000000",
	"0000000000000000000111111111111111111111111111100000000000000000",
	"0000000000000000011111111111111111111111111111111000000000000000",
	"0000000000000000111111111111111111111111111111111100000000000000",
	"0000000000000011111111111111111111111111111111111110000000000000",
	"0000000000000111111111111111111111111111111111111111000000000000",
	"0000000000001111111111111111111111111111111111111111100000000000",
	"0000000000011111111111111111111111111111111111111111110000000000",
	"0000000000111111111111111111111111111111111111111111111000000000",
	"0000000000111111111111111111111111111111111111111111111000000000",
	"0000000001111111111111111111111111111111111111111111111100000000",
	"0000000011111111111111111111111111111111111111111111111110000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000001111111111111111111111000000011111111111111111111111000000",
	"0000001111111111111111111100000000001111111111111111111111000000",
	"0000011111111111111111111000000000000011111111111111111111100000",
	"0000011111111111111111110000000000000001111111111111111111100000",
	"0000111111111111111111100000000000000001111111111111111111100000",
	"0000111111111111111111000000000000000000111111111111111111100000",
	"0000111111111111111110000000000000000000111111111111111111110000",
	"0001111111111111111110000000000000000000111111111111111111110000",
	"0001111111111111111110000000000000000000011111111111111111110000",
	"0001111111111111111100000000000000000000011111111111111000000000",
	"0011111111111111111100000000000000000000011111000000000000000000",
	"0011111111111111111100000000000000000000000000000000000000000000",
	"0011111111111111111000000000000000000000000000000000000000000000",
	"0011111111111111111000000000000000000000000000000000000000000000",
	"0011111111111111111000000000000000000000000000000000000000000000",
	"0111111111111111111000000000000000000000000000000000000000000000",
	"0111111111111111111000000000000000000000000000000000000000000000",
	"0111111111111111110000000000000000000000000000000000000000000000",
	"0111111111111111110000000000000000000000000000000000000000000000",
	"0111111111111111110000000000001111111111000000000000000000000000",
	"0111111111111111110000000011111111111111111000000000000000000000",
	"0111111111111111110000001111111111111111111111000000000000000000",
	"1111111111111111110000011111111111111111111111110000000000000000",
	"1111111111111111110001111111111111111111111111111000000000000000",
	"1111111111111111110011111111111111111111111111111100000000000000",
	"1111111111111111110111111111111111111111111111111111000000000000",
	"1111111111111111111111111111111111111111111111111111100000000000",
	"1111111111111111111111111111111111111111111111111111110000000000",
	"1111111111111111111111111111111111111111111111111111111000000000",
	"1111111111111111111111111111111111111111111111111111111000000000",
	"1111111111111111111111111111111111111111111111111111111100000000",
	"1111111111111111111111111111111111111111111111111111111110000000",
	"1111111111111111111111111111111111111111111111111111111111000000",
	"1111111111111111111111111111111111111111111111111111111111000000",
	"1111111111111111111111111111111111111111111111111111111111100000",
	"1111111111111111111111111110000000111111111111111111111111100000",
	"1111111111111111111111111000000000000111111111111111111111110000",
	"1111111111111111111111110000000000000011111111111111111111110000",
	"1111111111111111111111100000000000000001111111111111111111110000",
	"1111111111111111111111000000000000000000111111111111111111111000",
	"1111111111111111111110000000000000000000011111111111111111111000",
	"1111111111111111111110000000000000000000011111111111111111111000",
	"1111111111111111111100000000000000000000001111111111111111111000",
	"1111111111111111111100000000000000000000001111111111111111111100",
	"1111111111111111111100000000000000000000001111111111111111111100",
	"0111111111111111111000000000000000000000000111111111111111111100",
	"0111111111111111111000000000000000000000000111111111111111111100",
	"0111111111111111111000000000000000000000000111111111111111111100",
	"0111111111111111111000000000000000000000000111111111111111111100",
	"0111111111111111111000000000000000000000000111111111111111111100",
	"0111111111111111111000000000000000000000000111111111111111111100",
	"0111111111111111111000000000000000000000000111111111111111111100",
	"0011111111111111111000000000000000000000000111111111111111111100",
	"0011111111111111111000000000000000000000000111111111111111111100",
	"0011111111111111111000000000000000000000000111111111111111111100",
	"0011111111111111111100000000000000000000000111111111111111111100",
	"0011111111111111111100000000000000000000000111111111111111111100",
	"0001111111111111111100000000000000000000001111111111111111111000",
	"0001111111111111111110000000000000000000001111111111111111111000",
	"0001111111111111111110000000000000000000001111111111111111111000",
	"0000111111111111111111000000000000000000011111111111111111111000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000111111111111111111110000000000000000111111111111111111110000",
	"0000011111111111111111111000000000000001111111111111111111110000",
	"0000011111111111111111111100000000000111111111111111111111100000",
	"0000001111111111111111111111000000011111111111111111111111100000",
	"0000001111111111111111111111111111111111111111111111111111000000",
	"0000000111111111111111111111111111111111111111111111111111000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000000011111111111111111111111111111111111111111111111110000000",
	"0000000001111111111111111111111111111111111111111111111100000000",
	"0000000000111111111111111111111111111111111111111111111000000000",
	"0000000000011111111111111111111111111111111111111111110000000000",
	"0000000000001111111111111111111111111111111111111111100000000000",
	"0000000000000111111111111111111111111111111111111111000000000000",
	"0000000000000011111111111111111111111111111111111110000000000000",
	"0000000000000001111111111111111111111111111111111100000000000000",
	"0000000000000000111111111111111111111111111111111000000000000000",
	"0000000000000000001111111111111111111111111111100000000000000000",
	"0000000000000000000011111111111111111111111110000000000000000000",
	"0000000000000000000000011111111111111111110000000000000000000000",
	"0000000000000000000000000011111111111100000000000000000000000000");
	
	-- constante para matriz do n�mero 7
	constant valor7 : valor := (
	"0000000000000000000000000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000000000000000000000000",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111000",
	"1111111111111111111111111111111111111111111111111111111111111000",
	"1111111111111111111111111111111111111111111111111111111111110000",
	"1111111111111111111111111111111111111111111111111111111111100000",
	"1111111111111111111111111111111111111111111111111111111111000000",
	"0000000000000000000000000000000000000000011111111111111110000000",
	"0000000000000000000000000000000000000000111111111111111100000000",
	"0000000000000000000000000000000000000001111111111111111000000000",
	"0000000000000000000000000000000000000011111111111111111000000000",
	"0000000000000000000000000000000000000011111111111111110000000000",
	"0000000000000000000000000000000000000111111111111111100000000000",
	"0000000000000000000000000000000000001111111111111111100000000000",
	"0000000000000000000000000000000000011111111111111111000000000000",
	"0000000000000000000000000000000000011111111111111110000000000000",
	"0000000000000000000000000000000000111111111111111110000000000000",
	"0000000000000000000000000000000001111111111111111100000000000000",
	"0000000000000000000000000000000001111111111111111000000000000000",
	"0000000000000000000000000000000011111111111111111000000000000000",
	"0000000000000000000000000000000111111111111111110000000000000000",
	"0000000000000000000000000000000111111111111111110000000000000000",
	"0000000000000000000000000000001111111111111111100000000000000000",
	"0000000000000000000000000000001111111111111111000000000000000000",
	"0000000000000000000000000000011111111111111111000000000000000000",
	"0000000000000000000000000000111111111111111110000000000000000000",
	"0000000000000000000000000000111111111111111110000000000000000000",
	"0000000000000000000000000001111111111111111100000000000000000000",
	"0000000000000000000000000001111111111111111100000000000000000000",
	"0000000000000000000000000011111111111111111000000000000000000000",
	"0000000000000000000000000011111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111110000000000000000000000",
	"0000000000000000000000000111111111111111110000000000000000000000",
	"0000000000000000000000001111111111111111100000000000000000000000",
	"0000000000000000000000001111111111111111100000000000000000000000",
	"0000000000000000000000011111111111111111000000000000000000000000",
	"0000000000000000000000011111111111111111000000000000000000000000",
	"0000000000000000000000111111111111111111000000000000000000000000",
	"0000000000000000000000111111111111111110000000000000000000000000",
	"0000000000000000000000111111111111111110000000000000000000000000",
	"0000000000000000000001111111111111111100000000000000000000000000",
	"0000000000000000000001111111111111111100000000000000000000000000",
	"0000000000000000000011111111111111111100000000000000000000000000",
	"0000000000000000000011111111111111111000000000000000000000000000",
	"0000000000000000000011111111111111111000000000000000000000000000",
	"0000000000000000000111111111111111111000000000000000000000000000",
	"0000000000000000000111111111111111110000000000000000000000000000",
	"0000000000000000001111111111111111110000000000000000000000000000",
	"0000000000000000001111111111111111110000000000000000000000000000",
	"0000000000000000001111111111111111100000000000000000000000000000",
	"0000000000000000011111111111111111100000000000000000000000000000",
	"0000000000000000011111111111111111100000000000000000000000000000",
	"0000000000000000011111111111111111000000000000000000000000000000",
	"0000000000000000011111111111111111000000000000000000000000000000",
	"0000000000000000111111111111111111000000000000000000000000000000",
	"0000000000000000111111111111111111000000000000000000000000000000",
	"0000000000000000111111111111111110000000000000000000000000000000",
	"0000000000000001111111111111111110000000000000000000000000000000",
	"0000000000000001111111111111111110000000000000000000000000000000",
	"0000000000000001111111111111111110000000000000000000000000000000",
	"0000000000000001111111111111111100000000000000000000000000000000",
	"0000000000000001111111111111111100000000000000000000000000000000",
	"0000000000000011111111111111111100000000000000000000000000000000",
	"0000000000000011111111111111111100000000000000000000000000000000",
	"0000000000000011111111111111111100000000000000000000000000000000",
	"0000000000000011111111111111111100000000000000000000000000000000",
	"0000000000000011111111111111111000000000000000000000000000000000",
	"0000000000000111111111111111111000000000000000000000000000000000",
	"0000000000000111111111111111111000000000000000000000000000000000",
	"0000000000000111111111111111111000000000000000000000000000000000",
	"0000000000000111111111111111111000000000000000000000000000000000",
	"0000000000000111111111111111111000000000000000000000000000000000",
	"0000000000000111111111111111111000000000000000000000000000000000",
	"0000000000000111111111111111110000000000000000000000000000000000",
	"0000000000001111111111111111110000000000000000000000000000000000",
	"0000000000001111111111111111110000000000000000000000000000000000",
	"0000000000001111111111111111110000000000000000000000000000000000",
	"0000000000001111111111111111110000000000000000000000000000000000",
	"0000000000001111111111111111110000000000000000000000000000000000",
	"0000000000001111111111111111110000000000000000000000000000000000",
	"0000000000001111111111111111110000000000000000000000000000000000",
	"0000000000001111111111111111110000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000000000000000000000000");
	
	-- constante para matriz do n�mero 8
	constant valor8 : valor := (
	"0000000000000000000000000111111111111110000000000000000000000000",
	"0000000000000000000011111111111111111111111000000000000000000000",
	"0000000000000000001111111111111111111111111111000000000000000000",
	"0000000000000000111111111111111111111111111111110000000000000000",
	"0000000000000011111111111111111111111111111111111100000000000000",
	"0000000000001111111111111111111111111111111111111111000000000000",
	"0000000000011111111111111111111111111111111111111111100000000000",
	"0000000000111111111111111111111111111111111111111111110000000000",
	"0000000001111111111111111111111111111111111111111111111000000000",
	"0000000011111111111111111111111111111111111111111111111100000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000001111111111111111111111111111111111111111111111111111000000",
	"0000001111111111111111111111111111111111111111111111111111000000",
	"0000011111111111111111111111100000011111111111111111111111100000",
	"0000011111111111111111111110000000000111111111111111111111100000",
	"0000111111111111111111111000000000000001111111111111111111110000",
	"0000111111111111111111111000000000000000111111111111111111110000",
	"0000111111111111111111110000000000000000111111111111111111110000",
	"0001111111111111111111100000000000000000011111111111111111111000",
	"0001111111111111111111100000000000000000011111111111111111111000",
	"0001111111111111111111100000000000000000011111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0000111111111111111111000000000000000000001111111111111111110000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000011111111111111111100000000000000000011111111111111111100000",
	"0000011111111111111111110000000000000000111111111111111111100000",
	"0000011111111111111111110000000000000001111111111111111111000000",
	"0000001111111111111111111000000000000001111111111111111111000000",
	"0000000111111111111111111110000000000111111111111111111110000000",
	"0000000111111111111111111111100000011111111111111111111100000000",
	"0000000011111111111111111111111111111111111111111111111000000000",
	"0000000001111111111111111111111111111111111111111111110000000000",
	"0000000000111111111111111111111111111111111111111111100000000000",
	"0000000000001111111111111111111111111111111111111111000000000000",
	"0000000000000111111111111111111111111111111111111100000000000000",
	"0000000000000001111111111111111111111111111111111000000000000000",
	"0000000000000000001111111111111111111111111111000000000000000000",
	"0000000000000000111111111111111111111111111111110000000000000000",
	"0000000000000011111111111111111111111111111111111100000000000000",
	"0000000000001111111111111111111111111111111111111111000000000000",
	"0000000000011111111111111111111111111111111111111111100000000000",
	"0000000001111111111111111111111111111111111111111111111000000000",
	"0000000011111111111111111111111111111111111111111111111100000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000001111111111111111111111000000011111111111111111111111000000",
	"0000001111111111111111111100000000000011111111111111111111000000",
	"0000011111111111111111111000000000000001111111111111111111100000",
	"0000111111111111111111110000000000000000111111111111111111110000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0001111111111111111111100000000000000000011111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111110000000000000000000000111111111111111111110",
	"0111111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111111000000000000000000000111111111111111111100",
	"0011111111111111111111000000000000000000001111111111111111111100",
	"0011111111111111111111100000000000000000001111111111111111111000",
	"0001111111111111111111100000000000000000011111111111111111111000",
	"0001111111111111111111110000000000000000111111111111111111111000",
	"0000111111111111111111111000000000000001111111111111111111110000",
	"0000111111111111111111111110000000000011111111111111111111110000",
	"0000011111111111111111111111100000001111111111111111111111100000",
	"0000011111111111111111111111111111111111111111111111111111100000",
	"0000001111111111111111111111111111111111111111111111111111000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000000011111111111111111111111111111111111111111111111100000000",
	"0000000001111111111111111111111111111111111111111111111000000000",
	"0000000000111111111111111111111111111111111111111111110000000000",
	"0000000000001111111111111111111111111111111111111111100000000000",
	"0000000000000111111111111111111111111111111111111110000000000000",
	"0000000000000001111111111111111111111111111111111100000000000000",
	"0000000000000000111111111111111111111111111111110000000000000000",
	"0000000000000000000111111111111111111111111111000000000000000000",
	"0000000000000000000001111111111111111111111000000000000000000000",
	"0000000000000000000000000011111111111110000000000000000000000000");
	
	-- constante para matriz do n�mero 9
	constant valor9 : valor := (
	"0000000000000000000000001111111111100000000000000000000000000000",
	"0000000000000000000011111111111111111110000000000000000000000000",
	"0000000000000000011111111111111111111111110000000000000000000000",
	"0000000000000001111111111111111111111111111100000000000000000000",
	"0000000000000011111111111111111111111111111111000000000000000000",
	"0000000000001111111111111111111111111111111111100000000000000000",
	"0000000000011111111111111111111111111111111111110000000000000000",
	"0000000000111111111111111111111111111111111111111000000000000000",
	"0000000001111111111111111111111111111111111111111100000000000000",
	"0000000011111111111111111111111111111111111111111110000000000000",
	"0000000111111111111111111111111111111111111111111111000000000000",
	"0000001111111111111111111111111111111111111111111111100000000000",
	"0000011111111111111111111111111111111111111111111111110000000000",
	"0000011111111111111111111111111111111111111111111111111000000000",
	"0000111111111111111111111111111111111111111111111111111000000000",
	"0000111111111111111111111111111111111111111111111111111100000000",
	"0001111111111111111111111110000001111111111111111111111100000000",
	"0001111111111111111111111000000000001111111111111111111110000000",
	"0011111111111111111111110000000000000111111111111111111110000000",
	"0011111111111111111111100000000000000011111111111111111111000000",
	"0011111111111111111111000000000000000001111111111111111111000000",
	"0111111111111111111110000000000000000000111111111111111111000000",
	"0111111111111111111110000000000000000000111111111111111111100000",
	"0111111111111111111100000000000000000000011111111111111111100000",
	"0111111111111111111100000000000000000000011111111111111111100000",
	"1111111111111111111100000000000000000000001111111111111111110000",
	"1111111111111111111000000000000000000000001111111111111111110000",
	"1111111111111111111000000000000000000000001111111111111111110000",
	"1111111111111111111000000000000000000000000111111111111111110000",
	"1111111111111111111000000000000000000000000111111111111111110000",
	"1111111111111111111000000000000000000000000111111111111111111000",
	"1111111111111111111000000000000000000000000111111111111111111000",
	"1111111111111111111000000000000000000000000111111111111111111000",
	"1111111111111111111000000000000000000000000111111111111111111000",
	"1111111111111111111000000000000000000000000111111111111111111000",
	"1111111111111111111000000000000000000000000111111111111111111000",
	"1111111111111111111000000000000000000000000111111111111111111000",
	"1111111111111111111000000000000000000000000111111111111111111100",
	"1111111111111111111000000000000000000000000111111111111111111100",
	"0111111111111111111100000000000000000000000111111111111111111100",
	"0111111111111111111100000000000000000000001111111111111111111100",
	"0111111111111111111100000000000000000000001111111111111111111100",
	"0111111111111111111110000000000000000000001111111111111111111100",
	"0011111111111111111110000000000000000000011111111111111111111100",
	"0011111111111111111111000000000000000000011111111111111111111100",
	"0011111111111111111111000000000000000000111111111111111111111100",
	"0001111111111111111111100000000000000001111111111111111111111100",
	"0001111111111111111111110000000000000011111111111111111111111100",
	"0000111111111111111111111100000000000111111111111111111111111100",
	"0000111111111111111111111111000000111111111111111111111111111100",
	"0000011111111111111111111111111111111111111111111111111111111100",
	"0000001111111111111111111111111111111111111111111111111111111100",
	"0000001111111111111111111111111111111111111111111111111111111100",
	"0000000111111111111111111111111111111111111111111111111111111100",
	"0000000011111111111111111111111111111111111111111111111111111100",
	"0000000001111111111111111111111111111111111111111111111111111100",
	"0000000000111111111111111111111111111111111011111111111111111100",
	"0000000000001111111111111111111111111111110011111111111111111100",
	"0000000000000111111111111111111111111111100011111111111111111100",
	"0000000000000011111111111111111111111111000011111111111111111100",
	"0000000000000000111111111111111111111100000011111111111111111000",
	"0000000000000000000111111111111111110000000011111111111111111000",
	"0000000000000000000000111111111100000000000011111111111111111000",
	"0000000000000000000000000000000000000000000011111111111111111000",
	"0000000000000000000000000000000000000000000011111111111111111000",
	"0000000000000000000000000000000000000000000111111111111111111000",
	"0000000000000000000000000000000000000000000111111111111111111000",
	"0000000000000000000000000000000000000000000111111111111111110000",
	"0000000000000000000000000000000000000000000111111111111111110000",
	"0000000000000000000000000000000000000000000111111111111111110000",
	"0000000000000000000000000000000000000000001111111111111111110000",
	"0000000000000000111110000000000000000000001111111111111111110000",
	"0000000111111111111110000000000000000000001111111111111111100000",
	"0011111111111111111110000000000000000000011111111111111111100000",
	"0011111111111111111111000000000000000000011111111111111111100000",
	"0011111111111111111111000000000000000000011111111111111111000000",
	"0001111111111111111111000000000000000000111111111111111111000000",
	"0001111111111111111111100000000000000001111111111111111111000000",
	"0001111111111111111111100000000000000011111111111111111110000000",
	"0001111111111111111111110000000000000111111111111111111110000000",
	"0000111111111111111111111100000000001111111111111111111100000000",
	"0000111111111111111111111111000000111111111111111111111100000000",
	"0000111111111111111111111111111111111111111111111111111000000000",
	"0000011111111111111111111111111111111111111111111111111000000000",
	"0000011111111111111111111111111111111111111111111111110000000000",
	"0000001111111111111111111111111111111111111111111111100000000000",
	"0000001111111111111111111111111111111111111111111111000000000000",
	"0000000111111111111111111111111111111111111111111111000000000000",
	"0000000011111111111111111111111111111111111111111110000000000000",
	"0000000001111111111111111111111111111111111111111100000000000000",
	"0000000001111111111111111111111111111111111111111000000000000000",
	"0000000000111111111111111111111111111111111111100000000000000000",
	"0000000000011111111111111111111111111111111111000000000000000000",
	"0000000000000111111111111111111111111111111110000000000000000000",
	"0000000000000011111111111111111111111111111000000000000000000000",
	"0000000000000000111111111111111111111111100000000000000000000000",
	"0000000000000000001111111111111111111100000000000000000000000000",
	"0000000000000000000000111111111111000000000000000000000000000000");
	
	constant valorGG : valor := (
	"0000000000000000000000000011111111111100000000000000000000000000",
	"0000000000000000000000111111111111111111110000000000000000000000",
	"0000000000000000000011111111111111111111111100000000000000000000",
	"0000000000000000001111111111111111111111111111000000000000000000",
	"0000000000000000111111111111111111111111111111110000000000000000",
	"0000000000000001111111111111111111111111111111111000000000000000",
	"0000000000000111111111111111111111111111111111111100000000000000",
	"0000000000001111111111111111111111111111111111111111000000000000",
	"0000000000011111111111111111111111111111111111111111000000000000",
	"0000000000011111111111111111111111111111111111111111100000000000",
	"0000000000111111111111111111111111111111111111111111110000000000",
	"0000000001111111111111111111111111111111111111111111111000000000",
	"0000000001111111111111111111111111111111111111111111111000000000",
	"0000000011111111111111111111111111111111111111111111111100000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000001111111111111111111111100000011111111111111111111111000000",
	"0000001111111111111111111110000000000111111111111111111111000000",
	"0000001111111111111111111100000000000011111111111111111111000000",
	"0000011111111111111111111000000000000001111111111111111111100000",
	"0000011111111111111111110000000000000000111111111111111111100000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000111111111111111111000000000000000000001111111111111111110000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111110000000000000000000000111111111111111111000",
	"0001111111111111111110000000000000000000000111111111111111111000",
	"0001111111111111111110000000000000000000000111111111111111111000",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000001111111111111111111100",
	"0011111111111111111110000000000000000000011111111111111111111100",
	"0011111111111111111110000000000000000000111111111111111111111100",
	"0011111111111111111110000000000000000001111111111111111111111100",
	"0011111111111111111100000000000000000011111111111111111111111100",
	"0011111111111111111100000000000000000111111111111111111111111100",
	"0111111111111111111100000000000000001111111111111111111111111110",
	"0111111111111111111100000000000000011111111111111111111111111110",
	"0111111111111111111100000000000000111111111111111111111111111110",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0011111111111111111100000000000000000000000000000000000000000000",
	"0011111111111111111100000000001111111111111111111111111100000000",
	"0011111111111111111100000000001111111111111111111111111110000000",
	"0011111111111111111110000000001111111111111111111111111111000000",
	"0011111111111111111110000000001111111111111111111111111111100000",
	"0011111111111111111110000000001111111111111111111111111111110000",
	"0011111111111111111110000000011111111111111111111111111111110000",
	"0011111111111111111110000000011111111111111111111111111111110000",
	"0001111111111111111110000000111111111111111111111111111111110000",
	"0001111111111111111110000000111111111111111111111111111111110000",
	"0001111111111111111111000000111111111111111111111111111111110000",
	"0001111111111111111111000000111111111111111111111111111111110000",
	"0001111111111111111111000000111111111110000001111111111111110000",
	"0000111111111111111111100000011111111110000011101111111111110000",
	"0000111111111111111111100000111111111110000011111111111111110000",
	"0000111111111111111111100000011111111110000111111111111111110000",
	"0000011111111111111111110000000000000000000111111111111111110000",
	"0000011111111111111111111100000000000000000111111111111111110000",
	"0000011111111111111111111110000000000000000111111111111111100000",
	"0000001111111111111111111110000000000000000111111111111111000000",
	"0000001111111111111111111111100000000000000111111111111111000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000000011111111111111111111111111111111111111111111111100000000",
	"0000000011111111111111111111111111111111111111111111111000000000",
	"0000000001111111111111111111111111111111111111111111111000000000",
	"0000000000111111111111111111111111111111111111111111110000000000",
	"0000000000011111111111111111111111111111111111111111100000000000",
	"0000000000001111111111111111111111111111111111111111100000000000",
	"0000000000000111111111111111111111111111111111111111000000000000",
	"0000000000000011111111111111111111111111111111111110000000000000",
	"0000000000000001111111111111111111111111111111111000000000000000",
	"0000000000000000111111111111111111111111111111110000000000000000",
	"0000000000000000001111111111111111111111111111000000000000000000",
	"0000000000000000000011111111111111111111111100000000000000000000",
	"0000000000000000000000111111111111111111110000000000000000000000",
	"0000000000000000000000000011111111111100000000000000000000000000");


	constant valorLL : valor := (
	"0111111111111111111111111100000000000000000000000000000000000000",
	"0111111111111111111111111100000000000000000000000000000000000000",
	"0111111111111111111111111100000000000000000000000000000000000000",
	"0111111111111111111111111100000000000000000000000000000000000000",
	"0111111111111111111111111100000000000000000000000000000000000000",
	"0111111111111111111111111100000000000000000000000000000000000000",
	"0111111111111111111111111100000000000000000000000000000000000000",
	"0111111111111111111111111100000000000000000000000000000000000000",
	"0111111111111111111111111100000000000000000000000000000000000000",
	"0111111111111111111111111100000000000000000000000000000000000000",
	"0111111111111111111111111100000000000000000000000000000000000000",
	"0111111111111111111111111100000000000000000000000000000000000000",
	"0111111111111111111111111100000000000000000000000000000000000000",
	"0111111111111111111111111100000000000000000000000000000000000000",
	"0111111111111111111111111100000000000000000000000000000000000000",
	"0111111111111111111111111100000000000000000000000000000000000000",
	"0111111111111111111100000000000000000000000000000000000000000000",
	"0111111111111111100000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111000000000000000000000000000000000000000000000000",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110");
	
--constant color_num			: std_logic_vector (7 downto 0) :=("11100011");--3 bits para red,3 bits para gree,2 bits para blue
	
--	constant num					:integer:=10;

--	signal sorteio11			   : std_logic_vector(3 downto 0) ; -- armazera temporariamente o valor da dezena do primeiro valor sorteado
--	signal sorteio21				: std_logic_vector(3 downto 0) ; -- armazera temporariamente o valor da unidade do primeiro valor sorteado
--	signal sorteio31				: std_logic_vector(3 downto 0) ; -- armazera temporariamente o valor da dezena do segundo valor sorteado
--	signal sorteio41				: std_logic_vector(3 downto 0) ; -- armazera temporariamente o valor da unidade do segundo valor sorteado
--	signal sorteio51				: std_logic_vector(3 downto 0) ; -- armazera temporariamente o valor da dezena do terceiro valor sorteado
--	signal sorteio61				: std_logic_vector(3 downto 0) ; -- armazera temporariamente o valor da unidade do terceiro valor sorteado
--	signal sorteio12				: std_logic_vector(3 downto 0) ; -- armazera temporariamente o valor da dezena do quarto valor sorteado
--	signal sorteio22				: std_logic_vector(3 downto 0) ; -- armazera temporariamente o valor da unidade do quarto valor sorteado
--	signal sorteio32				: std_logic_vector(3 downto 0) ; -- armazera temporariamente o valor da dezena do quinto valor sorteado
--	signal sorteio42				: std_logic_vector(3 downto 0) ; -- armazera temporariamente o valor da unidade do quinto valor sorteado
--	signal sorteio52				: std_logic_vector(3 downto 0) ; -- armazera temporariamente o valor da dezena do sexto valor sorteado
--	signal sorteio62				: std_logic_vector(3 downto 0) ; -- armazera temporariamente o valor da unidade do sexto valor sorteado
	

--	signal quadrante : std_logic_vector(3 downto 0):="1111";
--	signal score : std_logic_vector(3 downto 0):="1110";  
	
	
	--configura��o para resolu��o 800x600
	--configura��o horizontal VGA 
		constant Harea				: integer :=800;
		constant Hfrontporch		: integer :=40;
		constant Hsyncpulse		: integer :=128;
		constant Hbackporch		: integer :=88;
		constant Hwholeline		: integer :=1056;
	--configura��o vertical VGA
		constant Varea				: integer :=600;
		constant Vfrontporch		: integer :=1;
		constant Vsyncpulse		: integer :=4;
		constant Vbackporch		: integer :=23;
		constant Vwholeline		: integer :=628;

		constant ajusteH 			: integer:= 216;
		constant ajusteV 			: integer:= 27;


begin
-- processo gerenciado pelo clock
process (clk) 
	variable horizontal_cont : integer :=0; -- variavel para mapeamento horizontal do VGA
	variable vertical_cont   : integer :=0; -- variavel para mapeamento vertical do VGA
	variable valor_mapa : valor; -- variavel responsavel por armazenar o mapa binario (dezena ou unidade) do numero sorteado
	variable valor_mapa_dezena : valor;
--	variable score : std_logic_vector(3 downto 0):="1110"; --(score)  variavel responsavel por armazenar o numero sorteado
begin
	if rising_edge(clk) then
		if (horizontal_cont >= Hsyncpulse+Hbackporch )
			and (horizontal_cont < Hsyncpulse+Hbackporch+Harea )
			and (vertical_cont >= Vsyncpulse+Vbackporch )
			and (vertical_cont < Vsyncpulse+Vbackporch+Varea )
			then
			--(onde X corresponde a um valor de 1 a 6 ou seis sorteios)
			--esse IF mapear� o espa�o onde cada n�mero ser� plotado
			--X de 1 a 6 (6 n�meros sorteados)
			--se a posi��o do sorteio for X o valor da dezena ou unidade sorteado ser� atribuido a variavel "sorteio(x,y)" 
			--o valor da dezena ou unidade sorteado � atribuido a variavel valor_sort  
			--onde a componente que gerencia os mapas binarios receber� esse valor
			--far� uma varredura na matriz binaria
			--se o valor do ponteiro de varredura for 1 ir� plotar um pixel da cor especificada, 
			--sen�o ir� plotar um pixel da cor de fundo
			if (vertical_cont>=250+ajusteV)
			and(vertical_cont<=348+ajusteV)
			and(horizontal_cont>=336+ajusteH)
			and(horizontal_cont<=464+ajusteH) then
			-- (x,y) = (1,1)	x= digito correspondente  y= posi��o correspondente
				
				--if(sorteio=1) then
			--		sorteio11<=dec;
			--	end if;
				
				--valor_sort:=sorteio11;
				
		--		if(sorteio>=1) then
					if(valor_mapa_dezena(vertical_cont-(250+ajusteV))(horizontal_cont-(336+ajusteH))='1') then
						red <= "110";--color_num(7 downto 5);
						green <= "110";--color_num(4 downto 2); -- cor do numero(dezena) (score)
						blue <= "00";--color_num(1 downto 0);
					elsif(valor_mapa(vertical_cont-(250+ajusteV))(horizontal_cont-(400+ajusteH))='1') then
						red <= "000";--color_num(7 downto 5);
						green <= "110";--color_num(4 downto 2); -- cor do numero(unidade) (score)
						blue <= "11";--color_num(1 downto 0);
					else 
						red <= "000";
						green <= "000";	-- cor de fundo do numero(para bits 0 da matriz)
						blue <= "00";
					end if;
		--		else
		--			red <= "111";--color_num(7 downto 5);
		--			green <="000";-- color_num(4 downto 2);
		--			blue <= "00";--color_num(1 downto 0);
		--		end if;
				
			elsif (vertical_cont>=0+ajusteV) -- ajuste segundo quadrante amarelo
						and(vertical_cont<=300+ajusteV)
						and(horizontal_cont>=0+ajusteH)
						and(horizontal_cont<=400+ajusteH)
						and(quadrante(1)='1') then
							red <= "111";
							green <= "111";
							blue <= "00";
			elsif (vertical_cont >= 300+ajusteV)--ajuste terceiro quadrante vermelho 
						and(vertical_cont<=600+ajusteV)
						and(horizontal_cont>=0+ajusteH)
						and(horizontal_cont<=400+ajusteH)
						and(quadrante(2)='1')then
							red <= "111";
							green <= "000";
							blue <= "00";
			elsif (vertical_cont >= 0+ajusteV)-- ajuste primeiro quadrante verde
						and(vertical_cont<=300+ajusteV)
						and(horizontal_cont>=400+ajusteH)
						and(horizontal_cont<=800+ajusteH)
						and(quadrante(0)='1') then
							red <= "000";
							green <= "111";
							blue <= "00";
			elsif (vertical_cont >= 300+ajusteV)-- ajuste quarto quadrante azul
						and(vertical_cont<=600+ajusteV)
						and(horizontal_cont>=400+ajusteH)
						and(horizontal_cont<=800+ajusteH)
						and(quadrante(3)='1')then
							red <= "000";
							green <= "100";
							blue <= "11";
							
			else
							 red<="000";
							 green<="000";
							 blue<="00";
			end if;
		else -- caso estiver fora da limita��o da tela
			red <= "000";
			green <= "000";
			blue <= "00";
		end if;
		--ir� gerar o pulso para sincronizar horizontalmente o VGA
		if (horizontal_cont > 0 )
		and (horizontal_cont < Hsyncpulse+1 )
		then
			hs <= '0';
		else
			hs <= '1';
		end if;
		--ir� gerar o pulso para sincronizar verticalmente o VGA
		if (vertical_cont > 0 ) 
		and (vertical_cont < Vsyncpulse+1 )
		then
			vs <= '0';
		else
			vs <= '1';
		end if;
		-- a cada pulso de sincroniza��o horizontal incrementa o contador de maperamento horizontal
		horizontal_cont := horizontal_cont+1; 
		
		if (horizontal_cont=Hwholeline) then
			-- a cada pulso de sincroniza��o vertical incrementa o contador de maperamento vertical
			vertical_cont := vertical_cont+1; 
			horizontal_cont := 0;
		end if;
		
		if (vertical_cont=Vwholeline) then
			vertical_cont := 0;
		end if;
	end if;
	-- mapeamentos binarios numericos
	-- valor_mapa recebe o valor correspondente do n�mero
	case scoreVGA is
		when 0 =>valor_mapa:=valor0; 
		when 1 =>valor_mapa:=valor1; 
		when 2 =>valor_mapa:=valor2; 
		when 3 =>valor_mapa:=valor3; 
		when 4 =>valor_mapa:=valor4; 
		when 5 =>valor_mapa:=valor5; 
		when 6 =>valor_mapa:=valor6; 
		when 7 =>valor_mapa:=valor7; 
		when 8 =>valor_mapa:=valor8; 
		when 9 =>valor_mapa:=valor9;
		when 10 =>valor_mapa:=valor0;
		when 11 =>valor_mapa:=valor1; 
		when 12 =>valor_mapa:=valor2; 
		when 13 =>valor_mapa:=valor3; 
		when 14 =>valor_mapa:=valor4;
		when 15 =>valor_mapa:=valorGG;
		when others =>valor_mapa:=valorLL;	
	end case;
	if (scoreVGA > 9 and scoreVGA < 15) then
		valor_mapa_dezena := valor1;
		elsif(scoreVGA < 10)then
		valor_mapa_dezena := valor0;
		elsif(scoreVGA = 15)then
		valor_mapa_dezena := valorGG;
		else
		valor_mapa_dezena :=valorLL;
	end if;
	
end process;

end Behavioral;
